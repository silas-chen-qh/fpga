module kry_filter(
    input   clk,
    input   rst_n
    input   key_in,
    output  reg key_flag,
    output  reg key_state
)

